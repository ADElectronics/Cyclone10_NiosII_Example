
module nios2 (
	clk_clk,
	gpio_export,
	reset_reset_n);	

	input		clk_clk;
	output	[3:0]	gpio_export;
	input		reset_reset_n;
endmodule
